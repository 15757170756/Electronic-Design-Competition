library verilog;
use verilog.vl_types.all;
entity FPGA_EP2C_vlg_tst is
end FPGA_EP2C_vlg_tst;
